module id(
    
);
endmodule