`define Stop 1'b1
`define NoStop 1'b0
`define ZeroWord 32'd0
`define ZeroBit 1'b0
