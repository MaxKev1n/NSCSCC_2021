`include "global_define.vh"
`timescale 1ns / 1ps
module mux4x32(
    input [31:0] a0,
    input [31:0] a1,
    input [31:0] a2,
    input [31:0] a3,
    input [1:0] s,
    output [31:0] res
);

    assign res = s == 2'b00 ? a0 : (s == 2'b01 ? a1 : (s == 2'b10 ? a2 : a3));

endmodule