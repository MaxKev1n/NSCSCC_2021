`define Stop 1'b1
`define NoStop 1'b0
`define ZeroWord 32'd0
`define ZeroBit 1'b0
`define ADDU  23'b10000000000000000000000
`define ADD   23'b01000000000000000000000
`define SUB   23'b00100000000000000000000
`define SUBU  23'b00010000000000000000000
`define AND   23'b00001000000000000000000
`define OR    23'b00000100000000000000000
`define XOR   23'b00000010000000000000000
`define NOR   23'b00000001000000000000000
`define SLT   23'b00000000100000000000000
`define SLTU  23'b00000000010000000000000
`define SLL   23'b00000000001000000000000
`define SRL   23'b00000000000100000000000
`define SRA   23'b00000000000010000000000
`define LUI   23'b00000000000001000000000
`define JUMP_BRANCH 23'b00000000000000100000000
`define MULT  23'b00000000000000010000000
`define MULTU 23'b00000000000000001000000
`define DIV   23'b00000000000000000100000
`define DIVU  23'b00000000000000000010000
`define MFHI  23'b00000000000000000001000
`define MFLO  23'b00000000000000000000100
`define MTHI  23'b00000000000000000000010
`define MTLO  23'b00000000000000000000001
`define MEM_LB  8'b10000000
`define MEM_LBU 8'b01000000
`define MEM_LH  8'b00100000
`define MEM_LHU 8'b00010000
`define MEM_LW  8'b00001000
`define MEM_SB  8'b00000100
`define MEM_SH  8'b00000010
`define MEM_SW  8'b00000001