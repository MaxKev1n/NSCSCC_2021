module mem(
    input clk,
    input reset,
    input [31:0] da,
    input [31:0] db,
    input write_mem,
    output [31:0] dout
);

    

endmodule