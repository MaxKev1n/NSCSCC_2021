module pc(
    input 
);
endmodule