module exe();
endmodule