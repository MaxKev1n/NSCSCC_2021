module ALU(
    input [14:0] ALUControl,
    input [31:0] da,
    input [31:0] db,

    output [31:0] dout
);
endmodule