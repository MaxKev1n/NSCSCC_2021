`define Stop 1'b1
`define NoStop 1'b0
`define ZeroWord 32'd0
`define ZeroBit 1'b0
`define ADDU 15'b100000000000000
`define ADD  15'b010000000000000
`define SUB  15'b001000000000000
`define SUBU 15'b000100000000000
`define AND  15'b000010000000000
`define OR   15'b000001000000000
`define XOR  15'b000000100000000
`define NOR  15'b000000010000000
`define SLT  15'b000000001000000
`define SLTU 15'b000000000100000
`define SLL  15'b000000000010000
`define SRL  15'b000000000001000
`define SRA  15'b000000000000100
`define LUI  15'b000000000000010
`define JUMP_BRANCH 15'b000000000000001